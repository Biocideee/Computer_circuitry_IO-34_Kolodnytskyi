library verilog;
use verilog.vl_types.all;
entity mux4to1 is
end mux4to1;
